module des(clk, in, reset, out);

   parameter WIDTH=8;
   
   input clk, in, reset;
   output [WIDTH-1:0] out;
   
   // Fill Here
endmodule
